module tb;
    initial begin
        run_test ("test");
    end
endmodule