package params_pkg;
parameter PROFUNDIDAD = 14;
endpackage
